package pa_gpu;


endpackage