module comb_multiplier_tb;

  logic [23:0] a;
  logic [23:0] b;
  logic [47:0] result;

  initial begin
    a = '1; // 6
    b = 24'b111111110000000011111111; // -4
    #10us;
    $display("%d(%b) * %d(%b) = %d(%b)", $signed(a), a, $signed(b), b, $signed(result), result);
    $stop;
  end


  comb_multiplier multiplier(
    .a(a),
    .b(b),
    .result(result)
  );

endmodule
